library verilog;
use verilog.vl_types.all;
entity template_vlg_tb is
end template_vlg_tb;
