module uart(clk);
endmodule
