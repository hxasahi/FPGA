library verilog;
use verilog.vl_types.all;
entity demo_vlg_tst is
end demo_vlg_tst;
