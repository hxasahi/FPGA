library verilog;
use verilog.vl_types.all;
entity demo_vlg_tb is
end demo_vlg_tb;
