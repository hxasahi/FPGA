module uart();
endmodule
