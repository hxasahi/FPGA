library verilog;
use verilog.vl_types.all;
entity uart_vlg_tb is
end uart_vlg_tb;
