library verilog;
use verilog.vl_types.all;
entity uart_vlg_tst is
end uart_vlg_tst;
